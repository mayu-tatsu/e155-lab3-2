module testbench_lab3_mt();

    

endmodule